----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:43:03 07/21/2015 
-- Design Name: 
-- Module Name:    fsmc_glue - A_fsmc_glue 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity fsmc2bram is
  Generic (
    BW : positive; -- block width
    BS : positive; -- block select
    DW : positive; -- data witdth
    AW : positive; -- total address width
    count : positive
  );
	Port (
    fsmc_clk : in std_logic; -- extenal clock generated by FSMC bus

    A : in STD_LOGIC_VECTOR (AW-1 downto 0);
    D : inout STD_LOGIC_VECTOR (DW-1 downto 0);
    NWE : in STD_LOGIC;
    NOE : in STD_LOGIC;
    NCE : in STD_LOGIC;
    NBL : in std_logic_vector (1 downto 0);

    bram_a   : out STD_LOGIC_VECTOR (count*BW-1 downto 0);
    bram_di  : in  STD_LOGIC_VECTOR (count*DW-1 downto 0);
    bram_do  : out STD_LOGIC_VECTOR (count*DW-1 downto 0);
    bram_en  : out STD_LOGIC_vector (count-1    downto 0);
    bram_we  : out std_logic_vector (count*2-1  downto 0);
    bram_clk : out std_logic_vector (count-1    downto 0)
  );
  
  function address2en(A : in std_logic_vector(AW-1 downto 0)) return std_logic_vector is
  begin
    return A(AW-1 downto BW);
  end address2en;
  
  function address2cnt(A : in std_logic_vector(AW-1 downto 0)) return std_logic_vector is
  begin
    return A(BW-1 downto 0);
  end address2cnt;

end fsmc2bram;

-------------------------
architecture beh of fsmc2bram is

type state_t is (IDLE, ADDR, WRITE1, READ1);
signal state : state_t := IDLE;

signal a_cnt : STD_LOGIC_VECTOR (BW-1 downto 0) := (others => '0');

signal do_common : STD_LOGIC_VECTOR (DW-1 downto 0) := (others => '0');
signal di_common : STD_LOGIC_VECTOR (DW-1 downto 0) := (others => '0');
signal we_common : STD_LOGIC_VECTOR (1 downto 0) := (others => '0');
signal en_common : STD_LOGIC := '0';
signal blk_select : STD_LOGIC_VECTOR (BS-1 downto 0);

begin

  fanout : for n in 0 to count-1 generate 
  begin
    bram_a  ((n+1)*BW-1 downto n*BW) <= a_cnt;
    bram_we ((n+1)*2-1  downto n*2)  <= we_common;
    bram_do ((n+1)*DW-1 downto n*DW) <= do_common;
  end generate;
  bram_clk <= (others => fsmc_clk);
  
  
  
  en_demux : entity work.demuxer
  generic map (
    AW => BS,
    DW => 1
  )
  PORT MAP (
    A    => blk_select,
    i(0) => en_common,
    o    => bram_en
  );



  di_mux : entity work.muxer
  generic map (
    AW => BS,
    DW => DW
  )
  PORT MAP (
    A => blk_select,
    i => bram_di,
    o => di_common
  );



  D <= di_common when (NCE = '0' and NOE = '0') else (others => 'Z');
  do_common <= D;
  
  
  
  process(fsmc_clk, NCE) begin
    if (NCE = '1') then
      en_common <= '0';
      we_common <= "00";
      state <= IDLE;
      
    elsif rising_edge(fsmc_clk) then
      case state is
      
      when IDLE =>
        if (NCE = '0') then 
          a_cnt <= address2cnt(A);
          blk_select <= address2en(A);
          state <= ADDR;
        end if;
        
      when ADDR =>
        if (NWE = '0') then
          state <= WRITE1;
        else
          state <= READ1;
          en_common <= '1';
          a_cnt <= a_cnt + 1;
        end if;

      when WRITE1 =>
        en_common <= '1';
        we_common <= not NBL;
        a_cnt <= a_cnt + 1;

      when READ1 =>
        a_cnt <= a_cnt + 1;

      end case;
    end if;
  end process;
end beh;




